// Copyright(C) 2020 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by an MIT license file distributed with this software package

module particle

pub struct Color {
mut:
	r byte
	g byte
	b byte
	a byte
}
